module cpu_module (
    input wire clk,
    input wire reset,
    output reg [31:0] data_out,
    output reg error_flag
);

// Internal signals
reg [31:0] internal_data;
reg [31:0] counter;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        data_out <= 32'b0;
        internal_data <= 32'b0;
        counter <= 32'b0;
        error_flag <= 1'b0;
    end else begin
        // Data output logic
        counter <= counter + 1;
        if (counter == 32'hFFFFFFFF) begin
            error_flag <= 1'b1; // Set error flag if counter overflows
        end else begin
            internal_data <= counter;
            data_out <= internal_data;
            error_flag <= 1'b0;
        end
    end
end

endmodule